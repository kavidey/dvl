`ifndef CONSTANTS
   `define CONSTANTS

    // H-Bridge States
    `define HB_HIGHZ 2'b00
    `define HB_DAMP  2'b01
    `define HB_OSCL  2'b10
`endif