package dvl_pkg;
      typedef enum logic [1:0] {HIGHZ, DAMP, OSCL} h_bridge_state_t;
endpackage